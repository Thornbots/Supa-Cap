** Profile: "SCHEMATIC1-PeePeePooPoo"  [ C:\Users\teaneyje\Documents\Supa-Cap\Design Files\Super Capacitor V1\Simulations\PSpice\SuperCap-CapBoard-PSpiceFiles\SCHEMATIC1\PeePeePooPoo.sim ] 

** Creating circuit file "PeePeePooPoo.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\teaneyje\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "C:\Users\teaneyje\OneDrive - Rose-Hulman Institute of Technology\Documents\Classes\RHIT_Libraries\Class.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 400 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
